// RoundingMode
`define RM_RNE  3'b000
`define RM_RTZ  3'b001
`define RM_RDN  3'b010
`define RM_RUP  3'b011
`define RM_RMM  3'b100
`define RM_DYN  3'b111